`include "uvm_pkg.sv"
import uvm_pkg::*;
`include "mealy_overlap_11010.v"
`include "mealy_overlap_11010_common.sv"
`include "mealy_overlap_11010_tx.sv"
`include "mealy_overlap_11010_intf.sv"
`include "mealy_overlap_11010_seq_lib.sv"
`include "mealy_overlap_11010_sqr.sv"
`include "mealy_overlap_11010_drv.sv"
`include "mealy_overlap_11010_mon.sv"
`include "mealy_overlap_11010_sub.sv"
`include "mealy_overlap_11010_agent.sv"
`include "mealy_overlap_11010_sbd.sv"
`include "mealy_overlap_11010_env.sv"
`include "test_lib.sv"
`include "top.sv"
