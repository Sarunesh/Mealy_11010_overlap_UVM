class base_seq extends uvm_sequence#(mealy_overlap_11010_tx);
	// Factory registration
	`uvm_object_utils(base_seq)

	// Constructor
	`NEW_OBJECT
endclass
