interface mealy_overlap_11010_intf(input reg clk, input reg rst);
	logic data_out;
	logic data_in;
endinterface
